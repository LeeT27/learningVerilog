

module cpu_tb;

    reg clk;
    reg reset;

    
    CPU cpu (
        .clk(clk),
        .reset(reset)
    );

    initial clk = 0;
    always #5 clk = ~clk;
    
    initial begin
        $dumpfile("wave.vcd");
        $dumpvars(0, cpu);

        reset = 1;
        #10;
        reset = 0;

        // Instructions
        cpu.f2.memory[0]  = 32'b000100_1000000_00001_00000000000000; // LOAD mem[64] -> R1
        cpu.f2.memory[1]  = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[2]  = 32'b000100_1000001_00001_00000000000000; // LOAD mem[65] -> R1
        cpu.f2.memory[3]  = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[4]  = 32'b000100_1000010_00001_00000000000000; // LOAD mem[66] -> R1
        cpu.f2.memory[5]  = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[6]  = 32'b000100_1000011_00001_00000000000000; // LOAD mem[67] -> R1
        cpu.f2.memory[7]  = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[8]  = 32'b000100_1000100_00001_00000000000000; // LOAD mem[68] -> R1
        cpu.f2.memory[9]  = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[10] = 32'b000100_1000101_00001_00000000000000; // LOAD mem[69] -> R1
        cpu.f2.memory[11] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[12] = 32'b000100_1000110_00001_00000000000000; // LOAD mem[70] -> R1
        cpu.f2.memory[13] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[14] = 32'b000100_1000111_00001_00000000000000; // LOAD mem[71] -> R1
        cpu.f2.memory[15] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[16] = 32'b000100_1001000_00001_00000000000000; // LOAD mem[72] -> R1
        cpu.f2.memory[17] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[18] = 32'b000100_1001001_00001_00000000000000; // LOAD mem[73] -> R1
        cpu.f2.memory[19] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[20] = 32'b000100_1001010_00001_00000000000000; // LOAD mem[74] -> R1
        cpu.f2.memory[21] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[22] = 32'b000100_1001011_00001_00000000000000; // LOAD mem[75] -> R1
        cpu.f2.memory[23] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[24] = 32'b000100_1001100_00001_00000000000000; // LOAD mem[76] -> R1
        cpu.f2.memory[25] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[26] = 32'b000100_1001101_00001_00000000000000; // LOAD mem[77] -> R1
        cpu.f2.memory[27] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[28] = 32'b000100_1001110_00001_00000000000000; // LOAD mem[78] -> R1
        cpu.f2.memory[29] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[30] = 32'b000100_1001111_00001_00000000000000; // LOAD mem[79] -> R1
        cpu.f2.memory[31] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[32] = 32'b000100_1010000_00001_00000000000000; // LOAD mem[80] -> R1
        cpu.f2.memory[33] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[34] = 32'b000100_1010001_00001_00000000000000; // LOAD mem[81] -> R1
        cpu.f2.memory[35] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[36] = 32'b000100_1010010_00001_00000000000000; // LOAD mem[82] -> R1
        cpu.f2.memory[37] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[38] = 32'b000100_1010011_00001_00000000000000; // LOAD mem[83] -> R1
        cpu.f2.memory[39] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[40] = 32'b000100_1010100_00001_00000000000000; // LOAD mem[84] -> R1
        cpu.f2.memory[41] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[42] = 32'b000100_1010101_00001_00000000000000; // LOAD mem[85] -> R1
        cpu.f2.memory[43] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[44] = 32'b000100_1010110_00001_00000000000000; // LOAD mem[86] -> R1
        cpu.f2.memory[45] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[46] = 32'b000100_1010111_00001_00000000000000; // LOAD mem[87] -> R1
        cpu.f2.memory[47] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[48] = 32'b000100_1011000_00001_00000000000000; // LOAD mem[88] -> R1
        cpu.f2.memory[49] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[50] = 32'b000100_1011001_00001_00000000000000; // LOAD mem[89] -> R1
        cpu.f2.memory[51] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2
        cpu.f2.memory[52] = 32'b000100_1011010_00001_00000000000000; // LOAD mem[90] -> R1
        cpu.f2.memory[53] = 32'b000000_00001_00010_00010_00000000000; // ADD R1 + R2 -> R2

        cpu.f2.memory[54] = 32'b000100_1011100_00011_00000000000000; // LOAD 60 -> R3
        cpu.f2.memory[55] = 32'b000100_1011101_00100_00000000000000; // LOAD 262 -> R4
        cpu.f2.memory[56] = 32'b000100_1011110_00101_00000000000000; // LOAD 10 -> R5

        cpu.f2.memory[57] = 32'b000010_00010_00101_00010_00000000000; // MULT R2 * R5 -> R2
        cpu.f2.memory[58] = 32'b000011_00010_00100_00010_00000000000; // DIV R2 / 262 -> R2

        cpu.f2.memory[59] = 32'b000011_00010_00011_00110_00000000000; // DIV R2 / R3 -> R6 minutes
        cpu.f2.memory[60] = 32'b000010_00110_00011_00111_00000000000; // MULT R6 * 60 -> R7 
        cpu.f2.memory[61] = 32'b000001_00010_00111_01000_00000000000; // SUB R2 - R7 -> R8
        cpu.f2.memory[62] = 32'b000101_1111110_00110_00000000000000; // STORE R6 -> memory[126]
        cpu.f2.memory[63] = 32'b000101_1111111_01000_00000000000000; // STORE R8 -> memory[127]
            

        // Data
        cpu.f2.memory[64]  = 32'b00000000000000000000000110100100; // 420
        cpu.f2.memory[65]  = 32'b00000000000000000000000110100111; // 423
        cpu.f2.memory[66]  = 32'b00000000000000000000000110100111; // 423
        cpu.f2.memory[67]  = 32'b00000000000000000000000111000000; // 448
        cpu.f2.memory[68]  = 32'b00000000000000000000000110111100; // 444
        cpu.f2.memory[69]  = 32'b00000000000000000000000110110010; // 434
        cpu.f2.memory[70]  = 32'b00000000000000000000000110101001; // 425
        cpu.f2.memory[71]  = 32'b00000000000000000000000111000000; // 448
        cpu.f2.memory[72]  = 32'b00000000000000000000000110110010; // 434
        cpu.f2.memory[73]  = 32'b00000000000000000000000110110000; // 432
        cpu.f2.memory[74]  = 32'b00000000000000000000000110101011; // 427
        cpu.f2.memory[75]  = 32'b00000000000000000000000110111011; // 443
        cpu.f2.memory[76]  = 32'b00000000000000000000000111000001; // 449
        cpu.f2.memory[77]  = 32'b00000000000000000000000110110001; // 433
        cpu.f2.memory[78]  = 32'b00000000000000000000000110100100; // 420
        cpu.f2.memory[79]  = 32'b00000000000000000000000110110011; // 435
        cpu.f2.memory[80]  = 32'b00000000000000000000000110111000; // 440
        cpu.f2.memory[81]  = 32'b00000000000000000000000110101010; // 428
        cpu.f2.memory[82]  = 32'b00000000000000000000000110111001; // 441
        cpu.f2.memory[83]  = 32'b00000000000000000000000110110011; // 435
        cpu.f2.memory[84]  = 32'b00000000000000000000000110100111; // 423
        cpu.f2.memory[85]  = 32'b00000000000000000000000110101010; // 426
        cpu.f2.memory[86]  = 32'b00000000000000000000000110110101; // 437
        cpu.f2.memory[87]  = 32'b00000000000000000000000110110100; // 436
        cpu.f2.memory[88]  = 32'b00000000000000000000000110100101; // 421
        cpu.f2.memory[89]  = 32'b00000000000000000000000110111011; // 443
        cpu.f2.memory[90]  = 32'b00000000000000000000000110101011; // 427
        cpu.f2.memory[91]  = 32'b00000000000000000000000000000000;
        cpu.f2.memory[92]  = 32'b00000000000000000000000000111100; //60
        cpu.f2.memory[93]  = 32'b00000000000000000000000100000110; //262
        cpu.f2.memory[94]  = 32'b00000000000000000000000000001010; //10
        cpu.f2.memory[95]  = 32'b00000000000000000000000000000000;
        cpu.f2.memory[96]  = 32'b00000000000000000000000000000000;
        cpu.f2.memory[97]  = 32'b00000000000000000000000000000000;
        cpu.f2.memory[98]  = 32'b00000000000000000000000000000000;
        cpu.f2.memory[99]  = 32'b00000000000000000000000000000000;
        cpu.f2.memory[100] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[101] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[102] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[103] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[104] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[105] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[106] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[107] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[108] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[109] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[110] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[111] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[112] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[113] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[114] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[115] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[116] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[117] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[118] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[119] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[120] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[121] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[122] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[123] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[124] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[125] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[126] = 32'b00000000000000000000000000000000;
        cpu.f2.memory[127] = 32'b00000000000000000000000000000000;
        #1000;

        $display("+---------------------------+");
        $display("|                           |");
        $display("|  Average mile time: %0d:%02d  |", cpu.f3.register[6], cpu.f2.memory[127]);
        $display("|                           |");
        $display("+---------------------------+");
        $stop;
    end



endmodule
